PK   �wU�
��  ��     cirkitFile.json�]�o��W
߫�"����]��[���&0h}��ک,��u��{I�q,��ǙI�M���G��3���e��_�͢�6��ת٭���-�泏�)?��o���a�Y���/�}�8���?'��URl?=l7զ]HY�vY�I��2�2/���ӄՂkQp��X�����gwg���]�K\��]���f��Y�DۼJ��U�t�����j���rjC��##�u���4I]�2�UQ'KV���u]��bK�q��sͨ�s$�S��#9C�1�1�+����$Ft���Yly��,j����M�R���OJ����(��A�i��U
��,82ge�XZ'UV��Sc�T�tg��Jmʚ#�I��#Ď\2H�(C�cV)u���%���m�|iM�U!u��ӪZ"����ȭ�#MG��B*G��r�~�i\8�@F�t�	�1�d�P�&P�CY�\���Jt�"
�?��g�\���p@I��E���L�uH�
��5Q� ������1rl� �����! ��1���(�=s`|����V�0CK�бMj�CǼd��Y�(� P�f(��Q�!�C�=��(��cP�6��4f�،�*̄�h��U�������3߱�LH"��刀9���7PY��?��=C���70�����0W�p��q��S{��	��,���U���Aޫ�}�v?���N�E�p�$\2.�s�J��"�hυ9�%��\���"��4�#/zY_Sf�64�e�k�eC�`�A�biZ�6�F��u�,À�Ѡ��i�l�l0��4(�G3�y�YS�żC1����Р�Q\k����_~�F)�44(�i�D��A�P4l�%��kO�6���W�7OO4�L���	M$pQ�hjx�!�fy��4a;m����i+N�NrpFtzw'7��\h�ryД㴍�f��MξSF�b�M�M�����t,͵M��6��h
lZ��l��AS�>4�D ���h��$�S�h�ڶ�&�6վm��<�s�$\	I�%#�H�h.��KN�:"�Ҡ�������� �� ��@��`�р�Ѡ�Ӡ��`sssssss"W�łłł��"���#<���'��\.b�<�s��p�υ/�8yD�:"�Ҡ���	OM�'��\.�8y��rQp�υF���'��\.^8y��B#���'��\�w��s��o��h�*�ݲ|>��j���am��\�6�mSV����J
�N���E���B̂D�Iu�����9`�V��f���B�w{sՑ#���!�#�?%�\	L�32��B��[�nϾ�����[�2�бU�y��f�\jl�M���T~226��De�^�O��/14���sD�02240|ĄX(c�h�Ϙ�����?�%M�i��L��(���8���0x	�q� Ù�S4����U���/6�!�2��$x��3oɦ�k�^x% #0�0�s" #A� ؀l\�r�c4�1��-��7R�&Z�P/:b&8����	D��ѓ"�J4�r�24�~9	��5^l�=)�kD��2����u�nyۦܯ6�����c}�/@߯Jl��Yx��ϑ���D�ϐ�}iO���l�z�E3f�	�s,�ұ<���ޮ�g �5eX8wU��";��l�XB	�Oc
`��c~(op�q��8G[h���XP�1�q�.�< j�α��cP�"��K�QYW�>�@T`l�q�,�"`�Q�&,ƻ*u��/�"��P}0Avc@�\p�zd��E�q"V\��g=�����D�+�t}�.�Հk�ak\�>`�u�v�m����E6x���_d����E�\�>PGD<p	�@�X���v��.����1pu�`�0OG�����0͂�as����lP�Rz�łk��E,2��>�A���a@��/|e�S�U��c����� .�"��C�O�7B~��������K�o=�E��hg�:��Mh��;u��lE�����{p߃�����=���}����=D'��!|�{����Z���]�b,�q ���b���G,��(<�'�?3v�զj=��g���L���W)�]	�ָ3 c��m�G�uj-Ǟ%�=	���S�z����8b½�w�cN�^��;j1�Qo�ĝ�[��!d�#I����Ƒ�V���@�Z4䑆q��{���8LŽ�y�a�У^Ɔ<1kq/�Gv�7S����B��*p�	���+aq�O>u�E��Z{�z`�}4������Š��ظ����I�ĸI��);6e�&ulR�&}l��&sl2��ؔ����l��t��t��=�O{�6��8#l<%�qJ�xN�㜰��Ia�Ya����p����b�T�\nm�ϝ���z�k=l+��*g��2�-�ish-9�V���x�PΞ,���+��X����� ���,����m���K���f�P5�����n�v/���H~��� �J���4;60�ٯ�w���B�Bn_�D�L
Q�$+J��%+�Җ�t���f��Mq��a�g�f�D��f�ꗏ���X5ź:^χ�1}#�9�Dz?��,֢қ��bt:���0~*��S�O �e@~
�� ��0~���i�'��2 ?�g`��*q-���g�̡�ˡ� �Cd$��@��p"�8D@q�, �Y �!� �Cd�B ��"�7D@o�, �Y �2���.�{����������6�a7�1×7&�93�&w>�����Ḯȳ�*��Ϙȓ�-e�;�yoZ1��{(�<�c��&���ʙ��Gw�Z�,֦x�MN���D�4��ĻuMl �T=�i�mݕG��D�����٧������Q��f����}c?�Ͼu>�ծ��S���oVΣ���v��������v��\�j~^�V�uu�����_5�b�5��Ov��m�����I�?��n����6���q���� �3*�L˹L���S~���U����-¬R�D�.�,�J�Rj���:�E��X�<�@���
S�3B���#�B���y�� :�s�y�	��g!��nu�L�#)��7O�8#;C��=^�/��Go���cK��}��&�L�"�R��VPͥ079�\4z܏�v����\�g���^Z��<1�M����Ȇ�ݨ�l�B��u�y���H%���u�g�%S�hǻ�LH�"U�9f�_���������fkKw9�K[�힩\;#*�Ϲ~�{������5���	��2uR�ie��g�`t��!�v+�w$�Yy���^h�(�5L<sќt��pN�67��f�EΜUO�e"�M�@׉R,�
k,3�P��"���1��R1��3ˢOٍr����r.Ru�r��-
�u�'g<4�%��L�v�);|�ۇ9��c�]6�v�7l����l?�u�,7��>V]"�v��M��]=�oÞ����z [|���O���Mն����>��?��oB_�fݣ8�f�w���� mӾ_mޕ]ӳ+::fզ�d,��x5��O��9~!�a�ڴ�m��c����n�s�?��}�Oݲ��oo?��]�	X��>���)�!2#�d]�u=�h���w��Rx��n�W�������LQ"�s@�6�8�M��v0:phb��H���g9N^r�d9=�3��'�I�Z���~l'�:'4	9��9�Iȟ��S�s���B�d*��E���I$��j�,l�R���+|4^!�ۢ��G7(��������tX+\�W��ү�J�_�S�L�C�J�6�3��]RA�Zj��р��G�����ӿ7zҦ�W�i�����(���[�I����S[�t�x��?M��:?*��A(�Px�=��8{/X�O�"A�"Z$(P�/�8S�|T�K�)�n��Έ�nH��H�vWEW�A����9���֩VE��g��#��:s�2��i���3%�گH�^#�ޟ�<���z��u�̯'2��#1�j"��Yۮ��? ����kd����C/S��O�Cֿ�C�
j�Z)�8�0Ra����UA��_�{ҧ��)�~�uC�dP+TךA��]��W9���,�u�+	���<;����a�JD��#���}�nP!���=ʇCP���������àJDP�r^���8�'ĨS%��b�ʕ���O���Xx�XP2 ����	�����Q�#���|9�a�*���^���Wa'���8�z�x�{�2��Y�8!�*\� ���j4b?ʈR,���=T�3��B4z��]���i�)`��2�T�����i]��˚N�Ա�ФJ'u�e��o«��(�UTo�a`O$��ŁC�+�����ue�4p/�#3a�!�wraT㚓#UϜ�*S�a��z�c��m�fe׻٭߮���oU�`7{��~��][}�����:��?PK
   �wU�
��  ��                   cirkitFile.jsonPK      =   �    